module Instruction_Memory(
  output reg[31 : 0] Instruction, 
  input[31: 0] Address
  );

  reg [31:0] data[0:100];

  
  initial begin
    data[0] = 32'b1110_00_1_1101_0_0000_0000_000000010100; //MOV 
    data[1] = 32'b1110_00_1_1101_0_0000_0001_101000000001; //MOV
    data[2] = 32'b1110_00_1_1101_0_0000_0010_000100000011; //MOV
    data[3] = 32'b1110_00_0_0100_1_0010_0011_000000000010; //ADDS
    data[4] = 32'b1110_00_0_0101_0_0000_0100_000000000000; //ADC
    data[5] = 32'b1110_00_0_0010_0_0100_0101_000100000100; //SUB
    data[6] = 32'b1110_00_0_0110_0_0000_0110_000010100000; //SBC
    data[7] = 32'b1110_00_0_1100_0_0101_0111_000101000010; //ORR
    data[8] = 32'b1110_00_0_0000_0_0111_1000_000000000011; //AND 
    data[9] = 32'b1110_00_0_1111_0_0000_1001_000000000110; //MVN 
    data[10] = 32'b1110_00_0_0001_0_0100_1010_000000000101; //EOR
    data[11] = 32'b1110_00_0_1010_1_1000_0000_000000000110; //CMP 
    data[12] = 32'b0001_00_0_0100_0_0001_0001_000000000001; //ADDNE
    data[13] = 32'b1110_00_0_1000_1_1001_0000_000000001000; //TST
    data[14] = 32'b0000_00_0_0100_0_0010_0010_000000000010; //ADDEQ
    data[15] = 32'b1110_00_1_1101_0_0000_0000_101100000001; //MOV
    data[16] = 32'b1110_01_0_0100_0_0000_0001_000000000000; //STR
    data[17] = 32'b1110_01_0_0100_1_0000_1011_000000000000; //LDR 
    data[18] = 32'b1110_01_0_0100_0_0000_0010_000000000100; //STR
    data[19] = 32'b1110_01_0_0100_0_0000_0011_000000001000; //STR
    data[20] = 32'b1110_01_0_0100_0_0000_0100_000000001101; //STR
    data[21] = 32'b1110_01_0_0100_0_0000_0101_000000010000; //STR
    data[22] = 32'b1110_01_0_0100_0_0000_0110_000000010100; //STR
    data[23] = 32'b1110_01_0_0100_1_0000_1010_000000000100; //LDR
    data[24] = 32'b1110_01_0_0100_0_0000_0111_000000011000; //STR
    data[25] = 32'b1110_00_1_1101_0_0000_0001_000000010000; //MOV Changed the value from 4 to 16 to observe the impact of cache.
    data[26] = 32'b1110_00_1_1101_0_0000_0010_000000000000; //MOV
    data[27] = 32'b1110_00_1_1101_0_0000_0011_000000000000; //MOV
    data[28] = 32'b1110_00_0_0100_0_0000_0100_000100000011; //ADD
    data[29] = 32'b1110_01_0_0100_1_0100_0101_000000000000; //LDR
    data[30] = 32'b1110_01_0_0100_1_0100_0110_000000000100; //LDR
    data[31] = 32'b1110_00_0_1010_1_0101_0000_000000000110; //CMP
    data[32] = 32'b1100_01_0_0100_0_0100_0110_000000000000; //STRGT
    data[33] = 32'b1100_01_0_0100_0_0100_0101_000000000100; //STRGT
    data[34] = 32'b1110_00_1_0100_0_0011_0011_000000000001; //ADD
    data[35] = 32'b1110_00_1_1010_1_0011_0000_000000000011; //CMP
    data[36] = 32'b1011_10_1_0_111111111111111111110111 ; //BLT
    data[37] = 32'b1110_00_1_0100_0_0010_0010_000000000001; //ADD
    data[38] = 32'b1110_00_0_1010_1_0010_0000_000000000001; //CMP
    data[39] = 32'b1011_10_1_0_111111111111111111110011 ; //BLT 
    data[40] = 32'b1110_01_0_0100_1_0000_0001_000000000000; //LDR
    data[41] = 32'b1110_01_0_0100_1_0000_0010_000000000100; //LDR
    data[42] = 32'b1110_01_0_0100_1_0000_0011_000000001000; //STR
    data[43] = 32'b1110_01_0_0100_1_0000_0100_000000001100; //STR
    data[44] = 32'b1110_01_0_0100_1_0000_0101_000000010000; //STR
    data[45] = 32'b1110_01_0_0100_1_0000_0110_000000010100; //STR
    data[46] = 32'b1110_10_1_0_111111111111111111111111 ; //B
  end

  always @(Address) begin
    Instruction = data[Address[31:2]];
  end

endmodule